
module pwm_system (
	clk_clk,
	pwm_gen_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	pwm_gen_0_external_connection_export;
	input		reset_reset_n;
endmodule
