
module my_system (
	clk_clk,
	custome_pio_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	custome_pio_0_external_connection_export;
	input		reset_reset_n;
endmodule
